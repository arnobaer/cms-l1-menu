-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_test_axo_v1_v3_v4

-- Unique ID of L1 Trigger Menu:
-- 9aa98d25-7a9a-42e5-94be-dd3cfddbdfa7

-- Unique ID of firmware implementation:
-- d0bd8481-ba3d-40b2-8d50-ae6beb21297c

-- Scale set:
-- scales_2024_05_15

-- VHDL producer
-- version: 2.20.0
-- hash value: 01d3461e956f1972cb9cbbbbb32745d60d52a3d208431bb6763622d65d6a8291

-- tmEventSetup
-- version: 0.13.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal axol1tl_trigger_i16 : std_logic;
    signal axol1tl_trigger_i18 : std_logic;
    signal axol1tl_trigger_i19 : std_logic;
    signal axol1tl_trigger_i8 : std_logic;

-- Signal definition for algorithms names
    signal l1_axo_loose_v1 : std_logic;
    signal l1_axo_tight_v1 : std_logic;
    signal l1_axo_v_tight_v1 : std_logic;
    signal l1_axo_tight : std_logic;

-- ========================================================